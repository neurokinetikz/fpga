//=============================================================================
// Coupling Susceptibility Module - v11.1a
//
// Computes coupling susceptibility chi(r) for frequency ratios using the
// Unified Boundary-Attractor Framework formula:
//
//   chi(r) = sum_{p,q coprime, q<=5} (1/q^2) * L(r - p/q, w_rational)
//          + sum_{n} w_phi * L(r - phi^n, w_phi)
//
// where L(x,w) = 1/(1 + (x/w)^2) is a Lorentzian with width w.
//
// Parameters:
//   - Farey depth: q <= 5 (55 fractions in range [0.5, 5.0])
//   - Lorentzian width (rational): w = 0.03
//   - Lorentzian width (phi): w = 0.05
//   - Phi weight: w_phi = 0.3
//   - Phi^n for n in [-2, 5]: 0.382, 0.618, 1.0, 1.618, 2.618, 4.236
//
// Key positions from computed LUT:
//   - Integer ratios (1, 2, 3, 4): HIGH chi ~0.77-0.98 -> BOUNDARIES
//   - Half-integer ratios (1.5, 2.5, 3.5): chi ~0.25-0.28 -> ATTRACTORS
//   - phi^0.5 = 1.272: chi = 0.134 -> ATTRACTOR (alpha band)
//   - phi^1.25 = 1.825: chi = 0.126 -> FALLBACK (most stable!)
//   - phi^1.5 = 2.058: chi = 0.270 (near 2:1 but escaped)
//   - 2:1 catastrophe (2.0): chi = 0.769 -> DANGER ZONE
//
// v11.0: Initial implementation with manually hardcoded LUT
// v11.1a: Systematic Farey fraction computation (55 rationals + 6 phi^n)
//=============================================================================
`timescale 1ns / 1ps

module coupling_susceptibility #(
    parameter WIDTH = 18,
    parameter FRAC = 14,
    parameter NUM_OSCILLATORS = 21,
    parameter ENABLE_ADAPTIVE = 1    // 0 = disabled (v10.5), 1 = enabled (v11.x)
)(
    input  wire clk,
    input  wire rst,
    input  wire clk_en,

    // Oscillator frequencies (OMEGA_DT values for each oscillator)
    // Packed: [20:0] where each is WIDTH bits
    input  wire signed [NUM_OSCILLATORS*WIDTH-1:0] omega_dt_packed,

    // Reference frequency for ratio computation (typically theta at ~152 OMEGA_DT)
    input  wire signed [WIDTH-1:0] omega_dt_reference,

    // Per-oscillator coupling susceptibility chi (Q14 format)
    // High chi = near integer ratio = unstable (boundary)
    // Low chi = near half-integer ratio = stable (attractor)
    output wire signed [NUM_OSCILLATORS*WIDTH-1:0] chi_packed,

    // Position classification for each oscillator
    // 00 = attractor (half-integer), 01 = boundary (integer),
    // 10 = quarter-integer fallback, 11 = other
    output wire [NUM_OSCILLATORS*2-1:0] position_class_packed,

    // Aggregate outputs
    output wire signed [WIDTH-1:0] chi_max,      // Maximum chi across all oscillators
    output wire signed [WIDTH-1:0] chi_min,      // Minimum chi (most stable)
    output wire [4:0] chi_max_index              // Which oscillator has max chi
);

//-----------------------------------------------------------------------------
// Constants
//-----------------------------------------------------------------------------
localparam signed [WIDTH-1:0] ONE_Q14 = 18'sd16384;
localparam signed [WIDTH-1:0] HALF_Q14 = 18'sd8192;

// Chi thresholds for classification (empirically tuned)
localparam signed [WIDTH-1:0] CHI_BOUNDARY_THRESH = 18'sd12288;  // 0.75 - boundary zone
localparam signed [WIDTH-1:0] CHI_ATTRACTOR_THRESH = 18'sd4096;  // 0.25 - attractor zone

// LUT parameters
// Index range: ratio from 0.5 to 4.0 in steps of 0.0125
// That's (4.0 - 0.5) / 0.0125 = 280 entries
// Index = (ratio_q14 - 8192) >> 5  (divide by 512 for step = 0.03125)
// Actually let's use coarser steps for efficiency: step = 1/64 = 0.015625
// Index = (ratio_q14 - 8192) >> 6  (256 entries for ratio 0.5 to 4.5)
localparam LUT_SIZE = 256;
localparam signed [WIDTH-1:0] RATIO_MIN = 18'sd8192;   // 0.5 in Q14
localparam signed [WIDTH-1:0] RATIO_MAX = 18'sd73728;  // 4.5 in Q14
localparam INDEX_SHIFT = 8;  // ratio_q14 >> 8 after offset

//-----------------------------------------------------------------------------
// Chi LUT - Farey Fraction Computed Values (v11.1a)
//
// Index i maps to ratio r = 0.5 + i/16 (step = 0.0625)
// chi(r) = sum_{p,q coprime, q<=5} (1/q^2) * L(r-p/q, 0.03)
//        + sum_n 0.3 * L(r - phi^n, 0.05)
//
// Farey fractions included (q <= 5, 55 total):
//   q=1: 1, 2, 3, 4, 5 (weight = 1.0)
//   q=2: 1/2, 3/2, 5/2, 7/2, 9/2, 11/2 (weight = 0.25)
//   q=3: 1/3, 2/3, 4/3, 5/3, ... (weight = 0.111)
//   q=4: 1/4, 3/4, 5/4, 7/4, ... (weight = 0.0625)
//   q=5: 1/5, 2/5, 3/5, 4/5, ... (weight = 0.04)
//
// Phi^n boundaries included (n = -2 to 5):
//   phi^-2=0.382, phi^-1=0.618, phi^0=1.0, phi^1=1.618
//   phi^2=2.618, phi^3=4.236
//-----------------------------------------------------------------------------

// Precomputed chi values (Q14 format)
// Generated by scripts/generate_chi_lut.py using:
//   chi(r) = sum_{p,q coprime, q<=5} (1/q^2) * L(r-p/q, 0.03)
//          + sum_n 0.3 * L(r - phi^n, 0.05)
// See scripts/chi_lut_values.vh for generation details.
reg signed [WIDTH-1:0] chi_lut [0:LUT_SIZE-1];

//-----------------------------------------------------------------------------
// LUT Initialization - v11.1a Farey Fraction Computed Values
//
// Key positions (ratio -> chi decimal):
//   1.0 (idx 32):  0.980 - INTEGER BOUNDARY (q=1)
//   2.0 (idx 96):  0.769 - 2:1 CATASTROPHE (q=1, most dangerous)
//   3.0 (idx 160): 0.768 - INTEGER BOUNDARY (q=1)
//   4.0 (idx 224): 0.773 - INTEGER BOUNDARY (q=1)
//   1.5 (idx 64):  0.281 - HALF-INT ATTRACTOR (q=2)
//   2.5 (idx 128): 0.279 - HALF-INT ATTRACTOR (q=2)
//   3.5 (idx 192): 0.247 - HALF-INT ATTRACTOR (q=2)
//   phi^0.5 = 1.272 (idx 49):  0.134 - ATTRACTOR (alpha band!)
//   phi^1.25 = 1.825 (idx 84): 0.126 - FALLBACK (most stable!)
//   phi^1 = 1.618 (idx 71):    0.326 - near 5/3 boundary
//   phi^1.5 = 2.058 (idx 99):  0.270 - escaped from 2:1
//   phi^2 = 2.618 (idx 135):   0.324 - between attractors
//   phi^2.5 = 3.330 (idx 181): 0.156 - ATTRACTOR
//-----------------------------------------------------------------------------
initial begin
    // Ratio 0.500 to 0.609 (indices 0-7)
    chi_lut[0] = 18'sd5063; chi_lut[1] = 18'sd4498; chi_lut[2] = 18'sd3762;
    chi_lut[3] = 18'sd3494; chi_lut[4] = 18'sd3651; chi_lut[5] = 18'sd4173;
    chi_lut[6] = 18'sd4932; chi_lut[7] = 18'sd5485;

    // Ratio 0.625 to 0.734 (indices 8-15) - near phi^-1 = 0.618
    chi_lut[8] = 18'sd5487; chi_lut[9] = 18'sd5127; chi_lut[10] = 18'sd4785;
    chi_lut[11] = 18'sd4286; chi_lut[12] = 18'sd3508; chi_lut[13] = 18'sd2941;
    chi_lut[14] = 18'sd2690; chi_lut[15] = 18'sd2691;

    // Ratio 0.750 to 0.859 (indices 16-23)
    chi_lut[16] = 18'sd2737; chi_lut[17] = 18'sd2571; chi_lut[18] = 18'sd2436;
    chi_lut[19] = 18'sd2412; chi_lut[20] = 18'sd2292; chi_lut[21] = 18'sd2152;
    chi_lut[22] = 18'sd2114; chi_lut[23] = 18'sd2174;

    // Ratio 0.875 to 0.984 (indices 24-31) - approaching 1.0 BOUNDARY
    chi_lut[24] = 18'sd2325; chi_lut[25] = 18'sd2580; chi_lut[26] = 18'sd2980;
    chi_lut[27] = 18'sd3606; chi_lut[28] = 18'sd4610; chi_lut[29] = 18'sd6279;
    chi_lut[30] = 18'sd9095; chi_lut[31] = 18'sd13292;

    // Ratio 1.000 to 1.109 (indices 32-39) - 1.0 INTEGER BOUNDARY
    chi_lut[32] = 18'sd16056; // 1.0 BOUNDARY - chi = 0.980
    chi_lut[33] = 18'sd13284; chi_lut[34] = 18'sd9078;
    chi_lut[35] = 18'sd6253; chi_lut[36] = 18'sd4575; chi_lut[37] = 18'sd3561;
    chi_lut[38] = 18'sd2924; chi_lut[39] = 18'sd2511;

    // Ratio 1.125 to 1.234 (indices 40-47)
    chi_lut[40] = 18'sd2241; chi_lut[41] = 18'sd2074; chi_lut[42] = 18'sd1993;
    chi_lut[43] = 18'sd2007; chi_lut[44] = 18'sd2118; chi_lut[45] = 18'sd2201;
    chi_lut[46] = 18'sd2179; chi_lut[47] = 18'sd2256;

    // Ratio 1.250 to 1.359 (indices 48-55) - phi^0.5 = 1.272 ATTRACTOR
    chi_lut[48] = 18'sd2344;
    chi_lut[49] = 18'sd2193; // phi^0.5 = 1.272 - chi = 0.134 ATTRACTOR
    chi_lut[50] = 18'sd2048; chi_lut[51] = 18'sd2096;
    chi_lut[52] = 18'sd2371; chi_lut[53] = 18'sd2728; chi_lut[54] = 18'sd2646;
    chi_lut[55] = 18'sd2300;

    // Ratio 1.375 to 1.484 (indices 56-63)
    chi_lut[56] = 18'sd2141; chi_lut[57] = 18'sd2175; chi_lut[58] = 18'sd2184;
    chi_lut[59] = 18'sd2112; chi_lut[60] = 18'sd2158; chi_lut[61] = 18'sd2408;
    chi_lut[62] = 18'sd2960; chi_lut[63] = 18'sd3894;

    // Ratio 1.500 to 1.609 (indices 64-71) - 3/2 HALF-INT + phi^1 BOUNDARY
    chi_lut[64] = 18'sd4602; // 1.5 = 3/2 ATTRACTOR - chi = 0.281
    chi_lut[65] = 18'sd4131; chi_lut[66] = 18'sd3464;
    chi_lut[67] = 18'sd3246; chi_lut[68] = 18'sd3441; chi_lut[69] = 18'sd3991;
    chi_lut[70] = 18'sd4771;
    chi_lut[71] = 18'sd5339; // phi^1 = 1.618 - chi = 0.326

    // Ratio 1.625 to 1.734 (indices 72-79)
    chi_lut[72] = 18'sd5353; chi_lut[73] = 18'sd5000; chi_lut[74] = 18'sd4663;
    chi_lut[75] = 18'sd4166; chi_lut[76] = 18'sd3387; chi_lut[77] = 18'sd2817;
    chi_lut[78] = 18'sd2561; chi_lut[79] = 18'sd2554;

    // Ratio 1.750 to 1.859 (indices 80-87) - phi^1.25 = 1.825 FALLBACK
    chi_lut[80] = 18'sd2589; chi_lut[81] = 18'sd2409; chi_lut[82] = 18'sd2254;
    chi_lut[83] = 18'sd2207;
    chi_lut[84] = 18'sd2057; // phi^1.25 = 1.825 - chi = 0.126 MOST STABLE!
    chi_lut[85] = 18'sd1878; chi_lut[86] = 18'sd1790; chi_lut[87] = 18'sd1785;

    // Ratio 1.875 to 1.984 (indices 88-95) - approaching 2:1 CATASTROPHE
    chi_lut[88] = 18'sd1848; chi_lut[89] = 18'sd1983; chi_lut[90] = 18'sd2216;
    chi_lut[91] = 18'sd2603; chi_lut[92] = 18'sd3262; chi_lut[93] = 18'sd4440;
    chi_lut[94] = 18'sd6610; chi_lut[95] = 18'sd10144;

    // Ratio 2.000 to 2.109 (indices 96-103) - 2:1 HARMONIC CATASTROPHE
    chi_lut[96] = 18'sd12600; // 2.0 = 2:1 CATASTROPHE - chi = 0.769
    chi_lut[97] = 18'sd10136; chi_lut[98] = 18'sd6594;
    chi_lut[99] = 18'sd4416; // phi^1.5 = 2.058 - chi = 0.270 (escaped!)
    chi_lut[100] = 18'sd3229; chi_lut[101] = 18'sd2560;
    chi_lut[102] = 18'sd2163; chi_lut[103] = 18'sd1918;

    // Ratio 2.125 to 2.234 (indices 104-111)
    chi_lut[104] = 18'sd1769; chi_lut[105] = 18'sd1690; chi_lut[106] = 18'sd1677;
    chi_lut[107] = 18'sd1742; chi_lut[108] = 18'sd1893; chi_lut[109] = 18'sd2008;
    chi_lut[110] = 18'sd2012; chi_lut[111] = 18'sd2110;

    // Ratio 2.250 to 2.359 (indices 112-119)
    chi_lut[112] = 18'sd2215; chi_lut[113] = 18'sd2079; chi_lut[114] = 18'sd1946;
    chi_lut[115] = 18'sd2004; chi_lut[116] = 18'sd2288; chi_lut[117] = 18'sd2653;
    chi_lut[118] = 18'sd2578; chi_lut[119] = 18'sd2237;

    // Ratio 2.375 to 2.484 (indices 120-127)
    chi_lut[120] = 18'sd2084; chi_lut[121] = 18'sd2122; chi_lut[122] = 18'sd2135;
    chi_lut[123] = 18'sd2067; chi_lut[124] = 18'sd2115; chi_lut[125] = 18'sd2369;
    chi_lut[126] = 18'sd2923; chi_lut[127] = 18'sd3860;

    // Ratio 2.500 to 2.609 (indices 128-135) - 5/2 HALF-INT + phi^2
    chi_lut[128] = 18'sd4569; // 2.5 = 5/2 ATTRACTOR - chi = 0.279
    chi_lut[129] = 18'sd4100; chi_lut[130] = 18'sd3434;
    chi_lut[131] = 18'sd3218; chi_lut[132] = 18'sd3414; chi_lut[133] = 18'sd3965;
    chi_lut[134] = 18'sd4746;
    chi_lut[135] = 18'sd5315; // phi^2 = 2.618 - chi = 0.324

    // Ratio 2.625 to 2.734 (indices 136-143)
    chi_lut[136] = 18'sd5330; chi_lut[137] = 18'sd4978; chi_lut[138] = 18'sd4642;
    chi_lut[139] = 18'sd4145; chi_lut[140] = 18'sd3367; chi_lut[141] = 18'sd2797;
    chi_lut[142] = 18'sd2541; chi_lut[143] = 18'sd2535;

    // Ratio 2.750 to 2.859 (indices 144-151)
    chi_lut[144] = 18'sd2570; chi_lut[145] = 18'sd2390; chi_lut[146] = 18'sd2235;
    chi_lut[147] = 18'sd2188; chi_lut[148] = 18'sd2038; chi_lut[149] = 18'sd1859;
    chi_lut[150] = 18'sd1771; chi_lut[151] = 18'sd1766;

    // Ratio 2.875 to 2.984 (indices 152-159) - approaching 3:1 BOUNDARY
    chi_lut[152] = 18'sd1829; chi_lut[153] = 18'sd1963; chi_lut[154] = 18'sd2196;
    chi_lut[155] = 18'sd2582; chi_lut[156] = 18'sd3241; chi_lut[157] = 18'sd4419;
    chi_lut[158] = 18'sd6588; chi_lut[159] = 18'sd10121;

    // Ratio 3.000 to 3.109 (indices 160-167) - 3:1 INTEGER BOUNDARY
    chi_lut[160] = 18'sd12577; // 3.0 BOUNDARY - chi = 0.768
    chi_lut[161] = 18'sd10112; chi_lut[162] = 18'sd6569;
    chi_lut[163] = 18'sd4390; chi_lut[164] = 18'sd3202; chi_lut[165] = 18'sd2531;
    chi_lut[166] = 18'sd2132; chi_lut[167] = 18'sd1886;

    // Ratio 3.125 to 3.234 (indices 168-175)
    chi_lut[168] = 18'sd1735; chi_lut[169] = 18'sd1654; chi_lut[170] = 18'sd1638;
    chi_lut[171] = 18'sd1701; chi_lut[172] = 18'sd1849; chi_lut[173] = 18'sd1961;
    chi_lut[174] = 18'sd1962; chi_lut[175] = 18'sd2055;

    // Ratio 3.250 to 3.359 (indices 176-183) - phi^2.5 = 3.330 ATTRACTOR
    chi_lut[176] = 18'sd2156; chi_lut[177] = 18'sd2015; chi_lut[178] = 18'sd1875;
    chi_lut[179] = 18'sd1927; chi_lut[180] = 18'sd2203;
    chi_lut[181] = 18'sd2558; // phi^2.5 = 3.330 - chi = 0.156 ATTRACTOR
    chi_lut[182] = 18'sd2472; chi_lut[183] = 18'sd2119;

    // Ratio 3.375 to 3.484 (indices 184-191)
    chi_lut[184] = 18'sd1949; chi_lut[185] = 18'sd1969; chi_lut[186] = 18'sd1959;
    chi_lut[187] = 18'sd1863; chi_lut[188] = 18'sd1877; chi_lut[189] = 18'sd2086;
    chi_lut[190] = 18'sd2583; chi_lut[191] = 18'sd3444;

    // Ratio 3.500 to 3.609 (indices 192-199) - 7/2 HALF-INT ATTRACTOR
    chi_lut[192] = 18'sd4053; // 3.5 = 7/2 ATTRACTOR - chi = 0.247
    chi_lut[193] = 18'sd3445; chi_lut[194] = 18'sd2583;
    chi_lut[195] = 18'sd2087; chi_lut[196] = 18'sd1878; chi_lut[197] = 18'sd1865;
    chi_lut[198] = 18'sd1961; chi_lut[199] = 18'sd1971;

    // Ratio 3.625 to 3.734 (indices 200-207)
    chi_lut[200] = 18'sd1952; chi_lut[201] = 18'sd2122; chi_lut[202] = 18'sd2476;
    chi_lut[203] = 18'sd2563; chi_lut[204] = 18'sd2208; chi_lut[205] = 18'sd1933;
    chi_lut[206] = 18'sd1882; chi_lut[207] = 18'sd2022;

    // Ratio 3.750 to 3.859 (indices 208-215)
    chi_lut[208] = 18'sd2165; chi_lut[209] = 18'sd2065; chi_lut[210] = 18'sd1973;
    chi_lut[211] = 18'sd1974; chi_lut[212] = 18'sd1864; chi_lut[213] = 18'sd1718;
    chi_lut[214] = 18'sd1657; chi_lut[215] = 18'sd1676;

    // Ratio 3.875 to 3.984 (indices 216-223) - approaching 4:1 BOUNDARY
    chi_lut[216] = 18'sd1760; chi_lut[217] = 18'sd1914; chi_lut[218] = 18'sd2164;
    chi_lut[219] = 18'sd2568; chi_lut[220] = 18'sd3244; chi_lut[221] = 18'sd4439;
    chi_lut[222] = 18'sd6627; chi_lut[223] = 18'sd10180;

    // Ratio 4.000 to 4.109 (indices 224-231) - 4:1 INTEGER BOUNDARY
    chi_lut[224] = 18'sd12658; // 4.0 BOUNDARY - chi = 0.773
    chi_lut[225] = 18'sd10218; chi_lut[226] = 18'sd6704;
    chi_lut[227] = 18'sd4559; chi_lut[228] = 18'sd3413; chi_lut[229] = 18'sd2796;
    chi_lut[230] = 18'sd2464; chi_lut[231] = 18'sd2306;

    // Ratio 4.125 to 4.234 (indices 232-239) - phi^3 = 4.236 BOUNDARY
    chi_lut[232] = 18'sd2274; chi_lut[233] = 18'sd2357; chi_lut[234] = 18'sd2572;
    chi_lut[235] = 18'sd2968; chi_lut[236] = 18'sd3591;
    chi_lut[237] = 18'sd4336; // near phi^3 = 4.236
    chi_lut[238] = 18'sd5014; chi_lut[239] = 18'sd5475;

    // Ratio 4.250 to 4.359 (indices 240-247)
    chi_lut[240] = 18'sd5332; chi_lut[241] = 18'sd4544; chi_lut[242] = 18'sd3746;
    chi_lut[243] = 18'sd3289; chi_lut[244] = 18'sd3206; chi_lut[245] = 18'sd3314;
    chi_lut[246] = 18'sd3053; chi_lut[247] = 18'sd2575;

    // Ratio 4.375 to 4.484 (indices 248-255)
    chi_lut[248] = 18'sd2314; chi_lut[249] = 18'sd2264; chi_lut[250] = 18'sd2202;
    chi_lut[251] = 18'sd2064; chi_lut[252] = 18'sd2045; chi_lut[253] = 18'sd2227;
    chi_lut[254] = 18'sd2702; chi_lut[255] = 18'sd3546;
end

//-----------------------------------------------------------------------------
// Unpack oscillator frequencies
//-----------------------------------------------------------------------------
wire signed [WIDTH-1:0] omega_dt [0:NUM_OSCILLATORS-1];
genvar g;
generate
    for (g = 0; g < NUM_OSCILLATORS; g = g + 1) begin : unpack_omega
        assign omega_dt[g] = omega_dt_packed[g*WIDTH +: WIDTH];
    end
endgenerate

//-----------------------------------------------------------------------------
// Per-oscillator chi computation
//-----------------------------------------------------------------------------
reg signed [WIDTH-1:0] chi_reg [0:NUM_OSCILLATORS-1];
reg [1:0] position_class_reg [0:NUM_OSCILLATORS-1];

// Ratio and LUT index computation
wire signed [2*WIDTH-1:0] ratio_full [0:NUM_OSCILLATORS-1];
wire signed [WIDTH-1:0] ratio_q14 [0:NUM_OSCILLATORS-1];
wire [7:0] lut_index [0:NUM_OSCILLATORS-1];
wire index_valid [0:NUM_OSCILLATORS-1];

generate
    for (g = 0; g < NUM_OSCILLATORS; g = g + 1) begin : ratio_calc
        // Ratio = omega_dt[g] / omega_dt_reference
        // For Q14 division: (omega_dt << 14) / reference
        assign ratio_full[g] = ({omega_dt[g], 14'b0}) /
                               (omega_dt_reference != 0 ? omega_dt_reference : 18'sd1);
        assign ratio_q14[g] = ratio_full[g][WIDTH-1:0];

        // LUT index: (ratio - 0.5) / 0.015625 = (ratio_q14 - 8192) >> 6
        // But we use >> 8 for 256 entries covering ratio 0.5 to 4.5
        wire signed [WIDTH-1:0] ratio_offset = ratio_q14[g] - RATIO_MIN;
        assign lut_index[g] = (ratio_offset[WIDTH-1]) ? 8'd0 :
                              (ratio_offset[WIDTH-1:INDEX_SHIFT] > 8'd255) ? 8'd255 :
                              ratio_offset[INDEX_SHIFT +: 8];
        assign index_valid[g] = (ratio_q14[g] >= RATIO_MIN) && (ratio_q14[g] <= RATIO_MAX);
    end
endgenerate

// Update chi values (registered for timing)
integer i;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        for (i = 0; i < NUM_OSCILLATORS; i = i + 1) begin
            chi_reg[i] <= 18'sd0;
            position_class_reg[i] <= 2'b11;  // Unknown
        end
    end else if (clk_en && ENABLE_ADAPTIVE) begin
        for (i = 0; i < NUM_OSCILLATORS; i = i + 1) begin
            // Read chi from LUT
            if (index_valid[i]) begin
                chi_reg[i] <= chi_lut[lut_index[i]];
            end else begin
                chi_reg[i] <= 18'sd8192;  // Default to 0.5 for out-of-range
            end

            // Classify position based on chi
            if (chi_reg[i] >= CHI_BOUNDARY_THRESH) begin
                position_class_reg[i] <= 2'b01;  // Boundary (integer)
            end else if (chi_reg[i] <= CHI_ATTRACTOR_THRESH) begin
                position_class_reg[i] <= 2'b00;  // Attractor (half-integer)
            end else if (chi_reg[i] <= 18'sd6554) begin
                position_class_reg[i] <= 2'b10;  // Quarter-integer fallback
            end else begin
                position_class_reg[i] <= 2'b11;  // Other
            end
        end
    end
end

//-----------------------------------------------------------------------------
// Pack outputs
//-----------------------------------------------------------------------------
generate
    for (g = 0; g < NUM_OSCILLATORS; g = g + 1) begin : pack_outputs
        assign chi_packed[g*WIDTH +: WIDTH] = ENABLE_ADAPTIVE ? chi_reg[g] : 18'sd0;
        assign position_class_packed[g*2 +: 2] = ENABLE_ADAPTIVE ? position_class_reg[g] : 2'b11;
    end
endgenerate

//-----------------------------------------------------------------------------
// Aggregate statistics
//-----------------------------------------------------------------------------
reg signed [WIDTH-1:0] chi_max_reg;
reg signed [WIDTH-1:0] chi_min_reg;
reg [4:0] chi_max_index_reg;

always @(posedge clk or posedge rst) begin
    if (rst) begin
        chi_max_reg <= 18'sd0;
        chi_min_reg <= ONE_Q14;
        chi_max_index_reg <= 5'd0;
    end else if (clk_en && ENABLE_ADAPTIVE) begin
        chi_max_reg <= 18'sd0;
        chi_min_reg <= ONE_Q14;
        chi_max_index_reg <= 5'd0;

        for (i = 0; i < NUM_OSCILLATORS; i = i + 1) begin
            if (chi_reg[i] > chi_max_reg) begin
                chi_max_reg <= chi_reg[i];
                chi_max_index_reg <= i[4:0];
            end
            if (chi_reg[i] < chi_min_reg) begin
                chi_min_reg <= chi_reg[i];
            end
        end
    end
end

assign chi_max = ENABLE_ADAPTIVE ? chi_max_reg : 18'sd0;
assign chi_min = ENABLE_ADAPTIVE ? chi_min_reg : 18'sd0;
assign chi_max_index = ENABLE_ADAPTIVE ? chi_max_index_reg : 5'd0;

endmodule
