//=============================================================================
// PV+ PING Network Testbench - v9.2
//
// Tests the Phase 3 PV+ interneuron model with dynamic state.
// Verifies:
// 1. PV+ state has temporal dynamics (leaky integrator)
// 2. PV+ phase lags pyramidal activity (~90 degrees)
// 3. E-I loop creates stable gamma oscillation
// 4. PV+ state resets properly
// 5. Comparison with expected tau = 5ms time constant
// 6. PING network behavior vs Phase 1 amplitude-proportional
//=============================================================================
`timescale 1ns / 1ps

module tb_pv_feedback;

parameter WIDTH = 18;
parameter FRAC = 14;
parameter FAST_SIM = 1;

reg clk;
reg rst;
reg clk_en;

// Cortical column inputs
reg signed [WIDTH-1:0] thalamic_theta_input;
reg signed [WIDTH-1:0] feedforward_input;
reg signed [WIDTH-1:0] matrix_thalamic_input;
reg signed [WIDTH-1:0] feedback_input_1;
reg signed [WIDTH-1:0] feedback_input_2;
reg signed [WIDTH-1:0] phase_couple_l23;
reg signed [WIDTH-1:0] phase_couple_l6;
reg encoding_window;
reg signed [WIDTH-1:0] mu_dt_l6, mu_dt_l5b, mu_dt_l5a, mu_dt_l4, mu_dt_l23;

// Cortical column outputs
wire signed [WIDTH-1:0] l23_x, l23_y;
wire signed [WIDTH-1:0] l5b_x, l5a_x;
wire signed [WIDTH-1:0] l6_x, l6_y;
wire signed [WIDTH-1:0] l4_x;

// Test tracking
integer test_num;
integer pass_count;
integer fail_count;
integer cycle_count;

// Amplitude tracking
reg signed [WIDTH-1:0] max_l23_amp;
reg signed [WIDTH-1:0] min_l23_amp;
wire signed [WIDTH-1:0] l23_amp;

// Compute amplitude approximation
wire signed [WIDTH-1:0] abs_x, abs_y;
assign abs_x = (l23_x < 0) ? -l23_x : l23_x;
assign abs_y = (l23_y < 0) ? -l23_y : l23_y;
assign l23_amp = (abs_x > abs_y) ? abs_x + (abs_y >>> 1) : abs_y + (abs_x >>> 1);

// Access internal PV+ state via hierarchical path
// v9.3: Signal renamed from pv_inhibition to pv_l23_inhibition
wire signed [WIDTH-1:0] pv_state;
wire signed [WIDTH-1:0] pv_inhibition;
assign pv_state = dut.pv_l23.pv_state;
assign pv_inhibition = dut.pv_l23_inhibition;

// Phase detection registers
reg signed [WIDTH-1:0] prev_l23_x;
reg signed [WIDTH-1:0] prev_pv_state;
integer l23_zero_cross_count;
integer pv_zero_cross_count;
integer l23_to_pv_phase_samples;
reg [31:0] phase_accumulator;

// Clock generation
initial begin
    clk = 0;
    forever #4 clk = ~clk;  // 125 MHz
end

// Clock enable generation
reg [3:0] clk_div;
always @(posedge clk) begin
    if (rst) begin
        clk_div <= 0;
        clk_en <= 0;
    end else begin
        clk_div <= clk_div + 1;
        clk_en <= (clk_div == 0);
    end
end

// DUT instantiation
cortical_column #(
    .WIDTH(WIDTH),
    .FRAC(FRAC)
) dut (
    .clk(clk),
    .rst(rst),
    .clk_en(clk_en),
    .thalamic_theta_input(thalamic_theta_input),
    .feedforward_input(feedforward_input),
    .matrix_thalamic_input(matrix_thalamic_input),
    .feedback_input_1(feedback_input_1),
    .feedback_input_2(feedback_input_2),
    .phase_couple_l23(phase_couple_l23),
    .phase_couple_l6(phase_couple_l6),
    .encoding_window(encoding_window),
    .attention_input(18'sd0),  // v9.4: No attention for PING tests
    .mu_dt_l6(mu_dt_l6),
    .mu_dt_l5b(mu_dt_l5b),
    .mu_dt_l5a(mu_dt_l5a),
    .mu_dt_l4(mu_dt_l4),
    .mu_dt_l23(mu_dt_l23),
    .l23_x(l23_x),
    .l23_y(l23_y),
    .l5b_x(l5b_x),
    .l5a_x(l5a_x),
    .l6_x(l6_x),
    .l6_y(l6_y),
    .l4_x(l4_x)
);

// Helper task: wait for N clk_en cycles
task wait_cycles;
    input integer n;
    integer i;
    begin
        for (i = 0; i < n; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);
        end
    end
endtask

// Helper task: run and track amplitude for N cycles
task run_and_track_amplitude;
    input integer n;
    integer i;
    begin
        max_l23_amp = 0;
        min_l23_amp = 18'sd32767;
        for (i = 0; i < n; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);
            if (l23_amp > max_l23_amp) max_l23_amp = l23_amp;
            if (l23_amp < min_l23_amp && l23_amp > 0) min_l23_amp = l23_amp;
        end
    end
endtask

// Helper task: count zero crossings
task count_zero_crossings;
    input integer n;
    integer i;
    begin
        l23_zero_cross_count = 0;
        pv_zero_cross_count = 0;
        prev_l23_x = l23_x;
        prev_pv_state = pv_state;

        for (i = 0; i < n; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);

            // Detect L2/3 zero crossing (positive going)
            if (prev_l23_x < 0 && l23_x >= 0) begin
                l23_zero_cross_count = l23_zero_cross_count + 1;
            end

            // Detect PV+ zero crossing (positive going)
            if (prev_pv_state < 0 && pv_state >= 0) begin
                pv_zero_cross_count = pv_zero_cross_count + 1;
            end

            prev_l23_x = l23_x;
            prev_pv_state = pv_state;
        end
    end
endtask

// Initialize inputs
task init_inputs;
    begin
        thalamic_theta_input = 0;
        feedforward_input = 0;
        matrix_thalamic_input = 0;
        feedback_input_1 = 0;
        feedback_input_2 = 0;
        phase_couple_l23 = 0;
        phase_couple_l6 = 0;
        encoding_window = 0;
        // Standard MU values
        mu_dt_l6 = 18'sd66;   // MU=4
        mu_dt_l5b = 18'sd66;
        mu_dt_l5a = 18'sd66;
        mu_dt_l4 = 18'sd66;
        mu_dt_l23 = 18'sd66;
    end
endtask

initial begin
    $display("=============================================================");
    $display("PV+ PING Network Testbench - v9.2");
    $display("=============================================================");

    test_num = 0;
    pass_count = 0;
    fail_count = 0;

    // Reset
    rst = 1;
    init_inputs;
    repeat(10) @(posedge clk);
    rst = 0;
    wait_cycles(10);

    //=========================================================================
    // Test 1: PV+ state resets to zero
    //=========================================================================
    test_num = 1;
    $display("\nTest %0d: PV+ state reset behavior", test_num);

    rst = 1;
    repeat(10) @(posedge clk);

    if (pv_state == 0) begin
        $display("  PASS: PV+ state resets to zero");
        pass_count = pass_count + 1;
    end else begin
        $display("  FAIL: PV+ state not zero after reset (got %0d)", pv_state);
        fail_count = fail_count + 1;
    end

    rst = 0;

    //=========================================================================
    // Test 2: PV+ state has dynamics (not instantaneous)
    //=========================================================================
    test_num = 2;
    $display("\nTest %0d: PV+ has temporal dynamics", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    feedforward_input = 18'sd4096;  // 0.25

    // Let system run briefly
    wait_cycles(50);

    begin : dynamics_test
        reg signed [WIDTH-1:0] pv_early;
        pv_early = pv_state;

        // Run more cycles
        wait_cycles(100);

        $display("  PV+ state early: %0d, later: %0d", pv_early, pv_state);

        // PV+ should change over time (dynamics)
        if (pv_state != pv_early) begin
            $display("  PASS: PV+ state evolves over time (has dynamics)");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: PV+ state static (no dynamics)");
            fail_count = fail_count + 1;
        end
    end

    //=========================================================================
    // Test 3: PV+ state varies dynamically (oscillation indicator)
    //=========================================================================
    test_num = 3;
    $display("\nTest %0d: PV+ state varies dynamically", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    feedforward_input = 18'sd4096;

    wait_cycles(500);  // Let oscillation stabilize

    // Track PV+ state variation over 500 cycles
    begin : pv_variation_test
        reg signed [WIDTH-1:0] pv_min, pv_max;
        integer i;

        pv_min = pv_state;
        pv_max = pv_state;

        for (i = 0; i < 500; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);
            if (pv_state < pv_min) pv_min = pv_state;
            if (pv_state > pv_max) pv_max = pv_state;
        end

        $display("  PV+ state range: min=%0d, max=%0d, span=%0d",
                 pv_min, pv_max, pv_max - pv_min);

        // PV+ has lowpass dynamics (tau=5ms), so it smooths gamma oscillation
        // Span > 100 indicates meaningful variation through the filter
        // The span is smaller than raw oscillation because of the filtering
        if ((pv_max - pv_min) > 100) begin
            $display("  PASS: PV+ state shows dynamic variation (filtered)");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: PV+ state too static");
            fail_count = fail_count + 1;
        end
    end

    //=========================================================================
    // Test 4: E-I loop creates stable gamma amplitude
    //=========================================================================
    test_num = 4;
    $display("\nTest %0d: E-I loop stabilizes gamma amplitude", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    feedforward_input = 18'sd4096;

    wait_cycles(500);

    run_and_track_amplitude(300);

    $display("  L2/3 amplitude range: min=%0d, max=%0d", min_l23_amp, max_l23_amp);

    // Amplitude should be bounded and stable
    if (max_l23_amp > 18'sd1000 && max_l23_amp < 18'sd35000) begin
        $display("  PASS: Gamma amplitude stable with PING network");
        pass_count = pass_count + 1;
    end else begin
        $display("  FAIL: Gamma amplitude not stable");
        fail_count = fail_count + 1;
    end

    //=========================================================================
    // Test 5: PV+ inhibition tracks pyramid output (with some delay)
    //=========================================================================
    test_num = 5;
    $display("\nTest %0d: PV+ tracks pyramid with temporal filtering", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    feedforward_input = 18'sd4096;

    wait_cycles(300);

    begin : tracking_test
        reg signed [WIDTH-1:0] l23_samples [0:9];  // Store last 10 pyramid samples
        reg signed [WIDTH-1:0] pv_sample;
        integer lag_correlation;
        integer instant_correlation;
        integer i, j;

        lag_correlation = 0;
        instant_correlation = 0;

        // Initialize sample buffer
        for (j = 0; j < 10; j = j + 1) l23_samples[j] = 0;

        // Sample relationship over multiple cycles
        for (i = 0; i < 100; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);

            // Shift sample buffer
            for (j = 9; j > 0; j = j - 1) l23_samples[j] = l23_samples[j-1];
            l23_samples[0] = l23_x;
            pv_sample = pv_state;

            // Instant correlation (same sign)
            if ((l23_samples[0] > 0 && pv_sample > 0) || (l23_samples[0] < 0 && pv_sample < 0))
                instant_correlation = instant_correlation + 1;

            // Lagged correlation (PV tracks where pyramid was 2 cycles ago)
            if (i >= 2) begin
                if ((l23_samples[2] > 0 && pv_sample > 0) || (l23_samples[2] < 0 && pv_sample < 0))
                    lag_correlation = lag_correlation + 1;
            end
        end

        $display("  Instant correlation: %0d/100, Lagged correlation: %0d/98",
                 instant_correlation, lag_correlation);

        // With tau=5ms at 4kHz update, response is relatively fast
        // PV should track pyramid closely (high correlation expected)
        // The key is that PV varies with pyramid, showing the feedback connection
        if (instant_correlation > 50) begin
            $display("  PASS: PV+ tracks pyramid activity");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: PV+ not tracking pyramid properly");
            fail_count = fail_count + 1;
        end
    end

    //=========================================================================
    // Test 6: High MU stability with PING network
    //=========================================================================
    test_num = 6;
    $display("\nTest %0d: High MU stability with PING", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    mu_dt_l23 = 18'sd99;  // MU=6 (high)
    feedforward_input = 18'sd4096;

    wait_cycles(500);

    run_and_track_amplitude(300);

    $display("  L2/3 amplitude with high MU: max=%0d", max_l23_amp);

    if (max_l23_amp < 18'sd45000) begin
        $display("  PASS: PING stabilizes high-MU oscillation");
        pass_count = pass_count + 1;
    end else begin
        $display("  FAIL: Amplitude too high with high MU");
        fail_count = fail_count + 1;
    end

    //=========================================================================
    // Test 7: Fast gamma (encoding window) with PING
    //=========================================================================
    test_num = 7;
    $display("\nTest %0d: Fast gamma stability with PING", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    encoding_window = 1;  // Fast gamma (65.3 Hz)
    feedforward_input = 18'sd4096;

    wait_cycles(500);

    run_and_track_amplitude(300);

    $display("  Fast gamma amplitude: max=%0d", max_l23_amp);

    if (max_l23_amp > 18'sd1000 && max_l23_amp < 18'sd35000) begin
        $display("  PASS: Fast gamma stable with PING network");
        pass_count = pass_count + 1;
    end else begin
        $display("  FAIL: Fast gamma not stable");
        fail_count = fail_count + 1;
    end

    //=========================================================================
    // Test 8: PV+ inhibition magnitude reasonable
    //=========================================================================
    test_num = 8;
    $display("\nTest %0d: PV+ inhibition magnitude", test_num);

    rst = 1;
    repeat(10) @(posedge clk);
    rst = 0;
    init_inputs;
    feedforward_input = 18'sd4096;

    wait_cycles(300);

    begin : inhibition_test
        reg signed [WIDTH-1:0] max_inhib;
        integer i;

        max_inhib = 0;
        for (i = 0; i < 200; i = i + 1) begin
            @(posedge clk);
            while (!clk_en) @(posedge clk);
            if (pv_inhibition > max_inhib) max_inhib = pv_inhibition;
            if (-pv_inhibition > max_inhib) max_inhib = -pv_inhibition;
        end

        $display("  Max PV+ inhibition: %0d", max_inhib);

        // Inhibition should be meaningful but not overwhelming
        if (max_inhib > 18'sd100 && max_inhib < 18'sd20000) begin
            $display("  PASS: PV+ inhibition in reasonable range");
            pass_count = pass_count + 1;
        end else begin
            $display("  FAIL: PV+ inhibition out of range");
            fail_count = fail_count + 1;
        end
    end

    //=========================================================================
    // Summary
    //=========================================================================
    $display("\n=============================================================");
    $display("PV+ PING Network Test Summary");
    $display("=============================================================");
    $display("Total tests: %0d", test_num);
    $display("Passed: %0d", pass_count);
    $display("Failed: %0d", fail_count);

    if (fail_count == 0) begin
        $display("\n*** ALL TESTS PASSED ***");
    end else begin
        $display("\n*** SOME TESTS FAILED ***");
    end

    $display("=============================================================");
    $finish;
end

endmodule
